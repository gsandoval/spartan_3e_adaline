----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Togno
-- 
-- Create Date:    18:45:51 07/05/2012 
-- Design Name: 
-- Module Name:    Adaline - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Adaline is
port(
	mclock : in std_logic;
	reset : in std_logic
);
end Adaline;

architecture Behavioral of Adaline is

begin


end Behavioral;

